/*
	��ɫ������ģ�飬����һ��ʱ�ӣ���������������Ƶĺ���ģʽ
*/
module tri_led (
	input wire clk,
	output wire tri_led0_r_n,	//��һ����ɫ�Ƶĺ�ɫ����
	output wire tri_led0_g_n,	//��һ����ɫ�Ƶ���ɫ����
	output wire tri_led0_b_n,	//��һ����ɫ�Ƶ���ɫ����
	output wire tri_led1_r_n,	//�ڶ�����ɫ�Ƶĺ�ɫ����
	output wire tri_led1_g_n,	//�ڶ�����ɫ�Ƶ���ɫ����
	output wire tri_led1_b_n	//�ڶ�����ɫ�Ƶ���ɫ����
);

endmodule
